module fetch

import net.http

fn fetch_pkgs() {
}
